module fulladder16 (A,B,SUM,CO);
	
	input [15:0]A;
	input [15:0]B;
	output CO;
	output [15:0]SUM;
	wire w1;
	wire w2;
	wire w3;

	rippleadd4bit c1( 1'b0, A[3:0], B[3:0], w1, SUM[3:0]);
	rippleadd4bit c2( w1, A[7:4], B[7:4], w2, SUM[7:4]);
	rippleadd4bit c3( w2, A[11:8], B[11:8], w3, SUM[11:8]);
	rippleadd4bit c4( w3, A[15:12], B[15:12], CO, SUM[15:12]);
   
endmodule 